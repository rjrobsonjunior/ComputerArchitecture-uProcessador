library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ULA_tb is
    port (
        clk   : in std_logic;
        reset : in std_logic;
        
    );
end entity;

architecture rtl of ULA_tb is

begin

    

end architecture;
