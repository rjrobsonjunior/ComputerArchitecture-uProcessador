library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
    port (
        clk     : in std_logic;
        address : in unsigned(6 downto 0);
        data    : out unsigned(15 downto 0)
    );
end entity;

architecture rtl of ROM is

    type mem is array (0 to 127) of unsigned(15  downto 0);
    constant rom_data : mem := (

    -- 0  => b"000000101_011_1000", -- ld r3, 5   (A)
    -- 1  => b"000001000_100_1000", -- ld r4, 8   (B)
    -- 2  => b"000000000_011_1101", -- movA r3    (C)
    -- 3  => b"000000000_100_0001", -- add r4     (C)
    -- 4  => b"000000000_101_1110", -- movR r5    (C)
    -- 5  => b"111111111_101_1001", -- addi -1    (D)
    -- 6  => b"000000000_101_1110", -- movR r5    (D)
    -- 7  => b"010100_000_000_1111", -- jump 0x14 (E)
    -- 8  => b"000000_000_101_1000", -- ld r5, 0  (F)
    -- 9  => x"F009", 
    -- 10  => x"F005",
    -- 11 => x"F007",
    -- 12  => x"9999",
    -- 13 => x"F000",
    -- 14 => x"0000",
    -- 15 => x"0000",
    -- 16 => x"0000",
    -- 17 => x"F009", 
    -- 18 => x"F005",
    -- 19 => x"F007",
    -- 20 => b"000000000_101_1101", -- movA r5    (G)
    -- 21 => b"000000000_011_1110", -- movR r3    (G)
    -- 22 => b"000010_000_011_1111", -- jump 0x02 (H)
    -- 23 => b"000000_000_101_1000", -- ld r5, 0  (I)

    -- 0  => b"000000000_011_1000", -- ld r3, 0   (A) x"0038"
    -- 1  => b"000000000_100_1000", -- ld r4, 0   (B) x"0048"
    -- 2  => b"000000000_011_1101", -- movA r3    (C) x"003D"
    -- 3  => b"000000000_100_0001", -- add r4     (C) x"0041"
    -- 4  => b"000000000_100_1110", -- movR r4    (D) x"003E"
    -- 5  => b"000000000_011_1101", -- movA r3    (D) x"003D"
    -- 6  => b"000000001_101_1001", -- addi 1     (D) x"00D9"
    -- 7  => b"000000000_011_1110", -- movR r3    (D) x"003E"
    -- 8  => b"000000011110_0111",  -- cmp 30     (E) x"01E7"
    -- 9  => b"111111111001_0101",  -- jz -7     (E) x"FD05"
    -- 10 => b"000000000_100_1101", -- movA r4    (F) x"004D"
    -- 11 => b"000000000_101_1110", -- movR r5    (F) x"005E"

    0  => b"001101001_001_1000", -- ld r1, 0x69
    1  => b"000000010_011_1000", -- ld r3, 2
    2  => b"000000000_001_1101", -- movA r1
    3  => b"000000000_011_1100", -- sw r3
    4  => b"000000000_000_1101", -- movA r0
    5  => b"000000000_011_1011", -- lw r3
    6  => b"000000000_000_1101", -- movA r0

    7  => b"000000001_111_1000", -- ld r7, 1
    8  => b"010101010_110_1000", -- ld r6, 0xAA
    9  => b"000000000_111_1101", -- movA r7
    10 => b"000000000_110_1100", -- sw r6
    11 => b"000000000_000_1101", -- movA r0
    12 => b"000000000_110_1011", -- lw r6
    13 => b"000000000_000_1101", -- movA r0

    14 => b"000001000_001_1000", -- ld r1, 8
    15 => b"000000000_000_1101", -- movA r0
    16 => b"010111010_000_1001", -- addi 0xBA
    17 => b"000000000_001_1100", -- sw r1
    18 => b"000000000_001_1101", -- movA r1
    19 => b"000000001_000_1101", -- addi 1
    20 => b"000000000_001_1110", -- movR r1

    21 => b"000001001_001_1000", -- ld r1, 9
    22 => b"000000000_000_1101", -- movA r0
    23 => b"010111010_000_1001", -- addi 0xBA
    24 => b"000000000_001_1100", -- sw r1
    25 => b"000000000_001_1101", -- movA r1
    26 => b"000000001_000_1101", -- addi 1
    27 => b"000000000_001_1110", -- movR r1

    28 => b"000001010_001_1000", -- ld r1, 10
    29 => b"000000000_000_1101", -- movA r0
    30 => b"011001010_000_1001", -- addi 0xCA
    31 => b"000000000_001_1100", -- sw r1

    32 => b"000001000_010_1000", -- ld r2, 8
    33 => b"000001001_011_1000", -- ld r3, 9
    34 => b"000001010_100_1000", -- ld r4, 10

    35 => b"000000000_010_1011", -- lw r2
    36 => b"000000000_000_1101", --movA r0

    37 => b"000000000_011_1011", -- lw r3
    38 => b"000000000_000_1101", --movA r0

    39 => b"000000000_100_1011", -- lw r4
    40 => b"000000000_000_1101", --movA r0
    others => (others => '0')
    );
begin
    process(clk)
    begin
        if(rising_edge(clk)) then
            data <= rom_data(to_integer(address));
        end if;
    end process;

end architecture;
